module top (
  input wire enable,
  input wire reset,
  input wire clk,
  output wire [127:0] O
);

wire [10:0] injector;


ro ro1 (
  .enable (enable),
  .inv (injector)
);

rg rg1 (
  .clk (clk),
  .enable (enable),
  .reset (reset),
  .injector (injector),
  .O (O)
);


endmodule


module ro (
  (*DONT_TOUCH= "true"*) input wire enable,
  (*DONT_TOUCH= "true"*) output wire O,
  (*DONT_TOUCH= "true"*) output wire[10:0] inv
);

  assign O = inv[0];

  (*DONT_TOUCH= "true"*) nand (inv[0], inv[1], enable);
  (*DONT_TOUCH= "true"*) not (inv[1], inv[2]);
  (*DONT_TOUCH= "true"*) not (inv[2], inv[3]);
  (*DONT_TOUCH= "true"*) not (inv[3], inv[4]);
  (*DONT_TOUCH= "true"*) not (inv[4], inv[5]);
  (*DONT_TOUCH= "true"*) not (inv[5], inv[6]);
  (*DONT_TOUCH= "true"*) not (inv[6], inv[7]);
  (*DONT_TOUCH= "true"*) not (inv[7], inv[8]);
  (*DONT_TOUCH= "true"*) not (inv[8], inv[9]);
  (*DONT_TOUCH= "true"*) not (inv[9], inv[10]);
  (*DONT_TOUCH= "true"*) not (inv[10], inv[0]);

endmodule


module rg (
  input wire clk,
  input wire enable,
  input wire reset,
  input wire [10:0] injector,
  output reg [255:0] O
);

wire example_internal_signal = 1'b0;

always @ (posedge clk or posedge reset) begin
  if (reset) begin
    O <= 256'd0;
  end else begin
    if (enable) begin
      O[0] <= O[1];
      O[1] <= O[2];
      O[2] <= O[3];
      O[3] <= O[4];
      O[4] <= O[5];
      O[5] <= O[6];
      O[6] <= O[7];
      O[7] <= O[8];
      O[8] <= O[9];
      O[9] <= O[10];
      O[10] <= O[11];
      O[11] <= O[12];
      O[12] <= O[13];
      O[13] <= O[14];
      O[14] <= O[15];
      O[15] <= O[16];
      O[16] <= O[17];
      O[17] <= O[18];
      O[18] <= O[19];
      O[19] <= O[20];
      O[20] <= O[21] ^ O[235];
      O[21] <= O[22];
      O[22] <= O[23];
      O[23] <= O[24];
      O[24] <= O[25];
      O[25] <= O[26];
      O[26] <= O[27];
      O[27] <= O[28];
      O[28] <= O[29];
      O[29] <= O[30];
      O[30] <= O[31];
      O[31] <= O[32];
      O[32] <= O[33];
      O[33] <= O[34];
      O[34] <= O[35];
      O[35] <= O[36];
      O[36] <= O[37];
      O[37] <= O[38];
      O[38] <= O[39];
      O[39] <= O[40];
      O[40] <= O[41];
      O[41] <= O[42];
      O[42] <= O[43] ^ O[213];
      O[43] <= O[44];
      O[44] <= O[45];
      O[45] <= O[46];
      O[46] <= O[47];
      O[47] <= O[48];
      O[48] <= O[49];
      O[49] <= O[50];
      O[50] <= O[51];
      O[51] <= O[52];
      O[52] <= O[53];
      O[53] <= O[54];
      O[54] <= O[55];
      O[55] <= O[56];
      O[56] <= O[57];
      O[57] <= O[58];
      O[58] <= O[59];
      O[59] <= O[60];
      O[60] <= O[61];
      O[61] <= O[62];
      O[62] <= O[63] ^ O[192];
      O[63] <= O[64];
      O[64] <= O[65];
      O[65] <= O[66];
      O[66] <= O[67];
      O[67] <= O[68];
      O[68] <= O[69];
      O[69] <= O[70];
      O[70] <= O[71];
      O[71] <= O[72];
      O[72] <= O[73];
      O[73] <= O[74];
      O[74] <= O[75];
      O[75] <= O[76];
      O[76] <= O[77];
      O[77] <= O[78];
      O[78] <= O[79];
      O[79] <= O[80];
      O[80] <= O[81];
      O[81] <= O[82];
      O[82] <= O[83];
      O[83] <= O[84] ^ O[171];
      O[84] <= O[85];
      O[85] <= O[86];
      O[86] <= O[87];
      O[87] <= O[88];
      O[88] <= O[89];
      O[89] <= O[90];
      O[90] <= O[91];
      O[91] <= O[92];
      O[92] <= O[93];
      O[93] <= O[94];
      O[94] <= O[95];
      O[95] <= O[96];
      O[96] <= O[97];
      O[97] <= O[98];
      O[98] <= O[99];
      O[99] <= O[100];
      O[100] <= O[101];
      O[101] <= O[102];
      O[102] <= O[103];
      O[103] <= O[104];
      O[104] <= O[105];
      O[105] <= O[106] ^ O[150];
      O[106] <= O[107];
      O[107] <= O[108];
      O[108] <= O[109];
      O[109] <= O[110];
      O[110] <= O[111];
      O[111] <= O[112];
      O[112] <= O[113];
      O[113] <= O[114];
      O[114] <= O[115];
      O[115] <= O[116];
      O[116] <= O[117];
      O[117] <= O[118];
      O[118] <= O[119];
      O[119] <= O[120];
      O[120] <= O[121];
      O[121] <= O[122];
      O[122] <= O[123];
      O[123] <= O[124];
      O[124] <= O[125];
      O[125] <= O[126];
      O[126] <= O[127];
      O[127] <= O[128];
      O[128] <= O[129];
      O[129] <= O[130];
      O[130] <= O[131];
      O[131] <= O[132];
      O[132] <= O[133];
      O[133] <= O[134];
      O[134] <= O[135];
      O[135] <= O[136];
      O[136] <= O[137];
      O[137] <= O[138];
      O[138] <= O[139];
      O[139] <= O[140];
      O[140] <= O[141];
      O[141] <= O[142];
      O[142] <= O[143];
      O[143] <= O[144];
      O[144] <= O[145];
      O[145] <= O[146];
      O[146] <= O[147];
      O[147] <= O[148];
      O[148] <= O[149];
      O[149] <= O[150];
      O[150] <= O[151];
      O[151] <= O[152];
      O[152] <= O[153];
      O[153] <= O[154];
      O[154] <= O[155];
      O[155] <= O[156];
      O[156] <= O[157];
      O[157] <= O[158];
      O[158] <= O[159];
      O[159] <= O[160];
      O[160] <= O[161];
      O[161] <= O[162];
      O[162] <= O[163];
      O[163] <= O[164];
      O[164] <= O[165];
      O[165] <= O[166];
      O[166] <= O[167];
      O[167] <= O[168];
      O[168] <= O[169];
      O[169] <= O[170];
      O[170] <= O[171];
      O[171] <= O[172];
      O[172] <= O[173];
      O[173] <= O[174];
      O[174] <= O[175];
      O[175] <= O[176];
      O[176] <= O[177];
      O[177] <= O[178];
      O[178] <= O[179];
      O[179] <= O[180];
      O[180] <= O[181];
      O[181] <= O[182];
      O[182] <= O[183];
      O[183] <= O[184];
      O[184] <= O[185];
      O[185] <= O[186];
      O[186] <= O[187];
      O[187] <= O[188];
      O[188] <= O[189];
      O[189] <= O[190];
      O[190] <= O[191];
      O[191] <= O[192];
      O[192] <= O[193];
      O[193] <= O[194];
      O[194] <= O[195];
      O[195] <= O[196];
      O[196] <= O[197];
      O[197] <= O[198];
      O[198] <= O[199];
      O[199] <= O[200];
      O[200] <= O[201];
      O[201] <= O[202];
      O[202] <= O[203];
      O[203] <= O[204];
      O[204] <= O[205];
      O[205] <= O[206];
      O[206] <= O[207];
      O[207] <= O[208];
      O[208] <= O[209];
      O[209] <= O[210];
      O[210] <= O[211];
      O[211] <= O[212];
      O[212] <= O[213];
      O[213] <= O[214];
      O[214] <= O[215];
      O[215] <= O[216];
      O[216] <= O[217];
      O[217] <= O[218];
      O[218] <= O[219];
      O[219] <= O[220];
      O[220] <= O[221];
      O[221] <= O[222];
      O[222] <= O[223];
      O[223] <= O[224];
      O[224] <= O[225];
      O[225] <= O[226];
      O[226] <= O[227];
      O[227] <= O[228];
      O[228] <= O[229];
      O[229] <= O[230];
      O[230] <= O[231];
      O[231] <= O[232];
      O[232] <= O[233];
      O[233] <= O[234];
      O[234] <= O[235];
      O[235] <= O[236];
      O[236] <= O[237];
      O[237] <= O[238];
      O[238] <= O[239];
      O[239] <= O[240];
      O[240] <= O[241];
      O[241] <= O[242];
      O[242] <= O[243];
      O[243] <= O[244];
      O[244] <= O[245] ^ injector[10];
      O[245] <= O[246] ^ injector[9];
      O[246] <= O[247] ^ injector[8];
      O[247] <= O[248] ^ injector[7];
      O[248] <= O[249] ^ injector[6];
      O[249] <= O[250] ^ injector[5];
      O[250] <= O[251] ^ injector[4];
      O[251] <= O[252] ^ injector[3];
      O[252] <= O[253] ^ injector[2];
      O[253] <= O[254] ^ injector[1];
      O[254] <= O[255] ^ injector[0];
      O[255] <= O[0];
    end
  end
end

endmodule