module tb (
);

  wire bist;
  wire clk_trng;
  wire enable;
  wire [255:0] injectors;
  wire [255:0] random_number;
  wire ready;
  wire reset;
  wire ro_clk;
  wire run;


  trng trng (
    .injectors ( injectors ),
    .rst ( reset ),
    .q ( random_number ),
    .clk ( clk_trng )
  );

  top fsm (
    .injectors ( injectors ),
    .reset ( reset ),
    .enable ( enable ),
    .ready ( ready ),
    .bist ( bist ),
    .run ( run ),
    .clk ( ro_clk )
  );

  clock_ro clock_ro (
    .en ( enable ),
    .clk ( ro_clk )
  );


  initial begin 
    $dumpfile("results/dump.vcd");
    $dumpvars(0,tb);
  end

  initial begin 
    #327690;
    $stop;
  end

  initial begin 
    force reset = 0;
    force bist = 0;
    force run = 0;
    #0.5;
    force reset = 1;
    #0.5;
    force reset = 0;
    force bist = 1;
    #0.5;
    force reset = 0;
    force run = 1;
    #0.5;
  end

// DFT_SIGNAL {injectors[0]}
// DFT_SIGNAL {injectors[1]}
// DFT_SIGNAL {injectors[2]}
// DFT_SIGNAL {injectors[3]}
// DFT_SIGNAL {injectors[4]}
// DFT_SIGNAL {injectors[5]}
// DFT_SIGNAL {injectors[6]}
// DFT_SIGNAL {injectors[7]}
// DFT_SIGNAL {injectors[8]}
// DFT_SIGNAL {injectors[9]}
// DFT_SIGNAL {injectors[10]}
// DFT_SIGNAL {injectors[11]}
// DFT_SIGNAL {injectors[12]}
// DFT_SIGNAL {injectors[13]}
// DFT_SIGNAL {injectors[14]}
// DFT_SIGNAL {injectors[15]}
// DFT_SIGNAL {injectors[16]}
// DFT_SIGNAL {injectors[17]}
// DFT_SIGNAL {injectors[18]}
// DFT_SIGNAL {injectors[19]}
// DFT_SIGNAL {injectors[20]}
// DFT_SIGNAL {injectors[21]}
// DFT_SIGNAL {injectors[22]}
// DFT_SIGNAL {injectors[23]}
// DFT_SIGNAL {injectors[24]}
// DFT_SIGNAL {injectors[25]}
// DFT_SIGNAL {injectors[26]}
// DFT_SIGNAL {injectors[27]}
// DFT_SIGNAL {injectors[28]}
// DFT_SIGNAL {injectors[29]}
// DFT_SIGNAL {injectors[30]}
// DFT_SIGNAL {injectors[31]}
// DFT_SIGNAL {injectors[32]}
// DFT_SIGNAL {injectors[33]}
// DFT_SIGNAL {injectors[34]}
// DFT_SIGNAL {injectors[35]}
// DFT_SIGNAL {injectors[36]}
// DFT_SIGNAL {injectors[37]}
// DFT_SIGNAL {injectors[38]}
// DFT_SIGNAL {injectors[39]}
// DFT_SIGNAL {injectors[40]}
// DFT_SIGNAL {injectors[41]}
// DFT_SIGNAL {injectors[42]}
// DFT_SIGNAL {injectors[43]}
// DFT_SIGNAL {injectors[44]}
// DFT_SIGNAL {injectors[45]}
// DFT_SIGNAL {injectors[46]}
// DFT_SIGNAL {injectors[47]}
// DFT_SIGNAL {injectors[48]}
// DFT_SIGNAL {injectors[49]}
// DFT_SIGNAL {injectors[50]}
// DFT_SIGNAL {injectors[51]}
// DFT_SIGNAL {injectors[52]}
// DFT_SIGNAL {injectors[53]}
// DFT_SIGNAL {injectors[54]}
// DFT_SIGNAL {injectors[55]}
// DFT_SIGNAL {injectors[56]}
// DFT_SIGNAL {injectors[57]}
// DFT_SIGNAL {injectors[58]}
// DFT_SIGNAL {injectors[59]}
// DFT_SIGNAL {injectors[60]}
// DFT_SIGNAL {injectors[61]}
// DFT_SIGNAL {injectors[62]}
// DFT_SIGNAL {injectors[63]}
// DFT_SIGNAL {injectors[64]}
// DFT_SIGNAL {injectors[65]}
// DFT_SIGNAL {injectors[66]}
// DFT_SIGNAL {injectors[67]}
// DFT_SIGNAL {injectors[68]}
// DFT_SIGNAL {injectors[69]}
// DFT_SIGNAL {injectors[70]}
// DFT_SIGNAL {injectors[71]}
// DFT_SIGNAL {injectors[72]}
// DFT_SIGNAL {injectors[73]}
// DFT_SIGNAL {injectors[74]}
// DFT_SIGNAL {injectors[75]}
// DFT_SIGNAL {injectors[76]}
// DFT_SIGNAL {injectors[77]}
// DFT_SIGNAL {injectors[78]}
// DFT_SIGNAL {injectors[79]}
// DFT_SIGNAL {injectors[80]}
// DFT_SIGNAL {injectors[81]}
// DFT_SIGNAL {injectors[82]}
// DFT_SIGNAL {injectors[83]}
// DFT_SIGNAL {injectors[84]}
// DFT_SIGNAL {injectors[85]}
// DFT_SIGNAL {injectors[86]}
// DFT_SIGNAL {injectors[87]}
// DFT_SIGNAL {injectors[88]}
// DFT_SIGNAL {injectors[89]}
// DFT_SIGNAL {injectors[90]}
// DFT_SIGNAL {injectors[91]}
// DFT_SIGNAL {injectors[92]}
// DFT_SIGNAL {injectors[93]}
// DFT_SIGNAL {injectors[94]}
// DFT_SIGNAL {injectors[95]}
// DFT_SIGNAL {injectors[96]}
// DFT_SIGNAL {injectors[97]}
// DFT_SIGNAL {injectors[98]}
// DFT_SIGNAL {injectors[99]}
// DFT_SIGNAL {injectors[100]}
// DFT_SIGNAL {injectors[101]}
// DFT_SIGNAL {injectors[102]}
// DFT_SIGNAL {injectors[103]}
// DFT_SIGNAL {injectors[104]}
// DFT_SIGNAL {injectors[105]}
// DFT_SIGNAL {injectors[106]}
// DFT_SIGNAL {injectors[107]}
// DFT_SIGNAL {injectors[108]}
// DFT_SIGNAL {injectors[109]}
// DFT_SIGNAL {injectors[110]}
// DFT_SIGNAL {injectors[111]}
// DFT_SIGNAL {injectors[112]}
// DFT_SIGNAL {injectors[113]}
// DFT_SIGNAL {injectors[114]}
// DFT_SIGNAL {injectors[115]}
// DFT_SIGNAL {injectors[116]}
// DFT_SIGNAL {injectors[117]}
// DFT_SIGNAL {injectors[118]}
// DFT_SIGNAL {injectors[119]}
// DFT_SIGNAL {injectors[120]}
// DFT_SIGNAL {injectors[121]}
// DFT_SIGNAL {injectors[122]}
// DFT_SIGNAL {injectors[123]}
// DFT_SIGNAL {injectors[124]}
// DFT_SIGNAL {injectors[125]}
// DFT_SIGNAL {injectors[126]}
// DFT_SIGNAL {injectors[127]}
// DFT_SIGNAL {injectors[128]}
// DFT_SIGNAL {injectors[129]}
// DFT_SIGNAL {injectors[130]}
// DFT_SIGNAL {injectors[131]}
// DFT_SIGNAL {injectors[132]}
// DFT_SIGNAL {injectors[133]}
// DFT_SIGNAL {injectors[134]}
// DFT_SIGNAL {injectors[135]}
// DFT_SIGNAL {injectors[136]}
// DFT_SIGNAL {injectors[137]}
// DFT_SIGNAL {injectors[138]}
// DFT_SIGNAL {injectors[139]}
// DFT_SIGNAL {injectors[140]}
// DFT_SIGNAL {injectors[141]}
// DFT_SIGNAL {injectors[142]}
// DFT_SIGNAL {injectors[143]}
// DFT_SIGNAL {injectors[144]}
// DFT_SIGNAL {injectors[145]}
// DFT_SIGNAL {injectors[146]}
// DFT_SIGNAL {injectors[147]}
// DFT_SIGNAL {injectors[148]}
// DFT_SIGNAL {injectors[149]}
// DFT_SIGNAL {injectors[150]}
// DFT_SIGNAL {injectors[151]}
// DFT_SIGNAL {injectors[152]}
// DFT_SIGNAL {injectors[153]}
// DFT_SIGNAL {injectors[154]}
// DFT_SIGNAL {injectors[155]}
// DFT_SIGNAL {injectors[156]}
// DFT_SIGNAL {injectors[157]}
// DFT_SIGNAL {injectors[158]}
// DFT_SIGNAL {injectors[159]}
// DFT_SIGNAL {injectors[160]}
// DFT_SIGNAL {injectors[161]}
// DFT_SIGNAL {injectors[162]}
// DFT_SIGNAL {injectors[163]}
// DFT_SIGNAL {injectors[164]}
// DFT_SIGNAL {injectors[165]}
// DFT_SIGNAL {injectors[166]}
// DFT_SIGNAL {injectors[167]}
// DFT_SIGNAL {injectors[168]}
// DFT_SIGNAL {injectors[169]}
// DFT_SIGNAL {injectors[170]}
// DFT_SIGNAL {injectors[171]}
// DFT_SIGNAL {injectors[172]}
// DFT_SIGNAL {injectors[173]}
// DFT_SIGNAL {injectors[174]}
// DFT_SIGNAL {injectors[175]}
// DFT_SIGNAL {injectors[176]}
// DFT_SIGNAL {injectors[177]}
// DFT_SIGNAL {injectors[178]}
// DFT_SIGNAL {injectors[179]}
// DFT_SIGNAL {injectors[180]}
// DFT_SIGNAL {injectors[181]}
// DFT_SIGNAL {injectors[182]}
// DFT_SIGNAL {injectors[183]}
// DFT_SIGNAL {injectors[184]}
// DFT_SIGNAL {injectors[185]}
// DFT_SIGNAL {injectors[186]}
// DFT_SIGNAL {injectors[187]}
// DFT_SIGNAL {injectors[188]}
// DFT_SIGNAL {injectors[189]}
// DFT_SIGNAL {injectors[190]}
// DFT_SIGNAL {injectors[191]}
// DFT_SIGNAL {injectors[192]}
// DFT_SIGNAL {injectors[193]}
// DFT_SIGNAL {injectors[194]}
// DFT_SIGNAL {injectors[195]}
// DFT_SIGNAL {injectors[196]}
// DFT_SIGNAL {injectors[197]}
// DFT_SIGNAL {injectors[198]}
// DFT_SIGNAL {injectors[199]}
// DFT_SIGNAL {injectors[200]}
// DFT_SIGNAL {injectors[201]}
// DFT_SIGNAL {injectors[202]}
// DFT_SIGNAL {injectors[203]}
// DFT_SIGNAL {injectors[204]}
// DFT_SIGNAL {injectors[205]}
// DFT_SIGNAL {injectors[206]}
// DFT_SIGNAL {injectors[207]}
// DFT_SIGNAL {injectors[208]}
// DFT_SIGNAL {injectors[209]}
// DFT_SIGNAL {injectors[210]}
// DFT_SIGNAL {injectors[211]}
// DFT_SIGNAL {injectors[212]}
// DFT_SIGNAL {injectors[213]}
// DFT_SIGNAL {injectors[214]}
// DFT_SIGNAL {injectors[215]}
// DFT_SIGNAL {injectors[216]}
// DFT_SIGNAL {injectors[217]}
// DFT_SIGNAL {injectors[218]}
// DFT_SIGNAL {injectors[219]}
// DFT_SIGNAL {injectors[220]}
// DFT_SIGNAL {injectors[221]}
// DFT_SIGNAL {injectors[222]}
// DFT_SIGNAL {injectors[223]}
// DFT_SIGNAL {injectors[224]}
// DFT_SIGNAL {injectors[225]}
// DFT_SIGNAL {injectors[226]}
// DFT_SIGNAL {injectors[227]}
// DFT_SIGNAL {injectors[228]}
// DFT_SIGNAL {injectors[229]}
// DFT_SIGNAL {injectors[230]}
// DFT_SIGNAL {injectors[231]}
// DFT_SIGNAL {injectors[232]}
// DFT_SIGNAL {injectors[233]}
// DFT_SIGNAL {injectors[234]}
// DFT_SIGNAL {injectors[235]}
// DFT_SIGNAL {injectors[236]}
// DFT_SIGNAL {injectors[237]}
// DFT_SIGNAL {injectors[238]}
// DFT_SIGNAL {injectors[239]}
// DFT_SIGNAL {injectors[240]}
// DFT_SIGNAL {injectors[241]}
// DFT_SIGNAL {injectors[242]}
// DFT_SIGNAL {injectors[243]}
// DFT_SIGNAL {injectors[244]}
// DFT_SIGNAL {injectors[245]}
// DFT_SIGNAL {injectors[246]}
// DFT_SIGNAL {injectors[247]}
// DFT_SIGNAL {injectors[248]}
// DFT_SIGNAL {injectors[249]}
// DFT_SIGNAL {injectors[250]}
// DFT_SIGNAL {injectors[251]}
// DFT_SIGNAL {injectors[252]}
// DFT_SIGNAL {injectors[253]}
// DFT_SIGNAL {injectors[254]}
// DFT_SIGNAL {injectors[255]}
// DFT_SIGNAL {reset}
// DFT_SIGNAL {random_number[0]}
// DFT_SIGNAL {random_number[1]}
// DFT_SIGNAL {random_number[2]}
// DFT_SIGNAL {random_number[3]}
// DFT_SIGNAL {random_number[4]}
// DFT_SIGNAL {random_number[5]}
// DFT_SIGNAL {random_number[6]}
// DFT_SIGNAL {random_number[7]}
// DFT_SIGNAL {random_number[8]}
// DFT_SIGNAL {random_number[9]}
// DFT_SIGNAL {random_number[10]}
// DFT_SIGNAL {random_number[11]}
// DFT_SIGNAL {random_number[12]}
// DFT_SIGNAL {random_number[13]}
// DFT_SIGNAL {random_number[14]}
// DFT_SIGNAL {random_number[15]}
// DFT_SIGNAL {random_number[16]}
// DFT_SIGNAL {random_number[17]}
// DFT_SIGNAL {random_number[18]}
// DFT_SIGNAL {random_number[19]}
// DFT_SIGNAL {random_number[20]}
// DFT_SIGNAL {random_number[21]}
// DFT_SIGNAL {random_number[22]}
// DFT_SIGNAL {random_number[23]}
// DFT_SIGNAL {random_number[24]}
// DFT_SIGNAL {random_number[25]}
// DFT_SIGNAL {random_number[26]}
// DFT_SIGNAL {random_number[27]}
// DFT_SIGNAL {random_number[28]}
// DFT_SIGNAL {random_number[29]}
// DFT_SIGNAL {random_number[30]}
// DFT_SIGNAL {random_number[31]}
// DFT_SIGNAL {random_number[32]}
// DFT_SIGNAL {random_number[33]}
// DFT_SIGNAL {random_number[34]}
// DFT_SIGNAL {random_number[35]}
// DFT_SIGNAL {random_number[36]}
// DFT_SIGNAL {random_number[37]}
// DFT_SIGNAL {random_number[38]}
// DFT_SIGNAL {random_number[39]}
// DFT_SIGNAL {random_number[40]}
// DFT_SIGNAL {random_number[41]}
// DFT_SIGNAL {random_number[42]}
// DFT_SIGNAL {random_number[43]}
// DFT_SIGNAL {random_number[44]}
// DFT_SIGNAL {random_number[45]}
// DFT_SIGNAL {random_number[46]}
// DFT_SIGNAL {random_number[47]}
// DFT_SIGNAL {random_number[48]}
// DFT_SIGNAL {random_number[49]}
// DFT_SIGNAL {random_number[50]}
// DFT_SIGNAL {random_number[51]}
// DFT_SIGNAL {random_number[52]}
// DFT_SIGNAL {random_number[53]}
// DFT_SIGNAL {random_number[54]}
// DFT_SIGNAL {random_number[55]}
// DFT_SIGNAL {random_number[56]}
// DFT_SIGNAL {random_number[57]}
// DFT_SIGNAL {random_number[58]}
// DFT_SIGNAL {random_number[59]}
// DFT_SIGNAL {random_number[60]}
// DFT_SIGNAL {random_number[61]}
// DFT_SIGNAL {random_number[62]}
// DFT_SIGNAL {random_number[63]}
// DFT_SIGNAL {random_number[64]}
// DFT_SIGNAL {random_number[65]}
// DFT_SIGNAL {random_number[66]}
// DFT_SIGNAL {random_number[67]}
// DFT_SIGNAL {random_number[68]}
// DFT_SIGNAL {random_number[69]}
// DFT_SIGNAL {random_number[70]}
// DFT_SIGNAL {random_number[71]}
// DFT_SIGNAL {random_number[72]}
// DFT_SIGNAL {random_number[73]}
// DFT_SIGNAL {random_number[74]}
// DFT_SIGNAL {random_number[75]}
// DFT_SIGNAL {random_number[76]}
// DFT_SIGNAL {random_number[77]}
// DFT_SIGNAL {random_number[78]}
// DFT_SIGNAL {random_number[79]}
// DFT_SIGNAL {random_number[80]}
// DFT_SIGNAL {random_number[81]}
// DFT_SIGNAL {random_number[82]}
// DFT_SIGNAL {random_number[83]}
// DFT_SIGNAL {random_number[84]}
// DFT_SIGNAL {random_number[85]}
// DFT_SIGNAL {random_number[86]}
// DFT_SIGNAL {random_number[87]}
// DFT_SIGNAL {random_number[88]}
// DFT_SIGNAL {random_number[89]}
// DFT_SIGNAL {random_number[90]}
// DFT_SIGNAL {random_number[91]}
// DFT_SIGNAL {random_number[92]}
// DFT_SIGNAL {random_number[93]}
// DFT_SIGNAL {random_number[94]}
// DFT_SIGNAL {random_number[95]}
// DFT_SIGNAL {random_number[96]}
// DFT_SIGNAL {random_number[97]}
// DFT_SIGNAL {random_number[98]}
// DFT_SIGNAL {random_number[99]}
// DFT_SIGNAL {random_number[100]}
// DFT_SIGNAL {random_number[101]}
// DFT_SIGNAL {random_number[102]}
// DFT_SIGNAL {random_number[103]}
// DFT_SIGNAL {random_number[104]}
// DFT_SIGNAL {random_number[105]}
// DFT_SIGNAL {random_number[106]}
// DFT_SIGNAL {random_number[107]}
// DFT_SIGNAL {random_number[108]}
// DFT_SIGNAL {random_number[109]}
// DFT_SIGNAL {random_number[110]}
// DFT_SIGNAL {random_number[111]}
// DFT_SIGNAL {random_number[112]}
// DFT_SIGNAL {random_number[113]}
// DFT_SIGNAL {random_number[114]}
// DFT_SIGNAL {random_number[115]}
// DFT_SIGNAL {random_number[116]}
// DFT_SIGNAL {random_number[117]}
// DFT_SIGNAL {random_number[118]}
// DFT_SIGNAL {random_number[119]}
// DFT_SIGNAL {random_number[120]}
// DFT_SIGNAL {random_number[121]}
// DFT_SIGNAL {random_number[122]}
// DFT_SIGNAL {random_number[123]}
// DFT_SIGNAL {random_number[124]}
// DFT_SIGNAL {random_number[125]}
// DFT_SIGNAL {random_number[126]}
// DFT_SIGNAL {random_number[127]}
// DFT_SIGNAL {random_number[128]}
// DFT_SIGNAL {random_number[129]}
// DFT_SIGNAL {random_number[130]}
// DFT_SIGNAL {random_number[131]}
// DFT_SIGNAL {random_number[132]}
// DFT_SIGNAL {random_number[133]}
// DFT_SIGNAL {random_number[134]}
// DFT_SIGNAL {random_number[135]}
// DFT_SIGNAL {random_number[136]}
// DFT_SIGNAL {random_number[137]}
// DFT_SIGNAL {random_number[138]}
// DFT_SIGNAL {random_number[139]}
// DFT_SIGNAL {random_number[140]}
// DFT_SIGNAL {random_number[141]}
// DFT_SIGNAL {random_number[142]}
// DFT_SIGNAL {random_number[143]}
// DFT_SIGNAL {random_number[144]}
// DFT_SIGNAL {random_number[145]}
// DFT_SIGNAL {random_number[146]}
// DFT_SIGNAL {random_number[147]}
// DFT_SIGNAL {random_number[148]}
// DFT_SIGNAL {random_number[149]}
// DFT_SIGNAL {random_number[150]}
// DFT_SIGNAL {random_number[151]}
// DFT_SIGNAL {random_number[152]}
// DFT_SIGNAL {random_number[153]}
// DFT_SIGNAL {random_number[154]}
// DFT_SIGNAL {random_number[155]}
// DFT_SIGNAL {random_number[156]}
// DFT_SIGNAL {random_number[157]}
// DFT_SIGNAL {random_number[158]}
// DFT_SIGNAL {random_number[159]}
// DFT_SIGNAL {random_number[160]}
// DFT_SIGNAL {random_number[161]}
// DFT_SIGNAL {random_number[162]}
// DFT_SIGNAL {random_number[163]}
// DFT_SIGNAL {random_number[164]}
// DFT_SIGNAL {random_number[165]}
// DFT_SIGNAL {random_number[166]}
// DFT_SIGNAL {random_number[167]}
// DFT_SIGNAL {random_number[168]}
// DFT_SIGNAL {random_number[169]}
// DFT_SIGNAL {random_number[170]}
// DFT_SIGNAL {random_number[171]}
// DFT_SIGNAL {random_number[172]}
// DFT_SIGNAL {random_number[173]}
// DFT_SIGNAL {random_number[174]}
// DFT_SIGNAL {random_number[175]}
// DFT_SIGNAL {random_number[176]}
// DFT_SIGNAL {random_number[177]}
// DFT_SIGNAL {random_number[178]}
// DFT_SIGNAL {random_number[179]}
// DFT_SIGNAL {random_number[180]}
// DFT_SIGNAL {random_number[181]}
// DFT_SIGNAL {random_number[182]}
// DFT_SIGNAL {random_number[183]}
// DFT_SIGNAL {random_number[184]}
// DFT_SIGNAL {random_number[185]}
// DFT_SIGNAL {random_number[186]}
// DFT_SIGNAL {random_number[187]}
// DFT_SIGNAL {random_number[188]}
// DFT_SIGNAL {random_number[189]}
// DFT_SIGNAL {random_number[190]}
// DFT_SIGNAL {random_number[191]}
// DFT_SIGNAL {random_number[192]}
// DFT_SIGNAL {random_number[193]}
// DFT_SIGNAL {random_number[194]}
// DFT_SIGNAL {random_number[195]}
// DFT_SIGNAL {random_number[196]}
// DFT_SIGNAL {random_number[197]}
// DFT_SIGNAL {random_number[198]}
// DFT_SIGNAL {random_number[199]}
// DFT_SIGNAL {random_number[200]}
// DFT_SIGNAL {random_number[201]}
// DFT_SIGNAL {random_number[202]}
// DFT_SIGNAL {random_number[203]}
// DFT_SIGNAL {random_number[204]}
// DFT_SIGNAL {random_number[205]}
// DFT_SIGNAL {random_number[206]}
// DFT_SIGNAL {random_number[207]}
// DFT_SIGNAL {random_number[208]}
// DFT_SIGNAL {random_number[209]}
// DFT_SIGNAL {random_number[210]}
// DFT_SIGNAL {random_number[211]}
// DFT_SIGNAL {random_number[212]}
// DFT_SIGNAL {random_number[213]}
// DFT_SIGNAL {random_number[214]}
// DFT_SIGNAL {random_number[215]}
// DFT_SIGNAL {random_number[216]}
// DFT_SIGNAL {random_number[217]}
// DFT_SIGNAL {random_number[218]}
// DFT_SIGNAL {random_number[219]}
// DFT_SIGNAL {random_number[220]}
// DFT_SIGNAL {random_number[221]}
// DFT_SIGNAL {random_number[222]}
// DFT_SIGNAL {random_number[223]}
// DFT_SIGNAL {random_number[224]}
// DFT_SIGNAL {random_number[225]}
// DFT_SIGNAL {random_number[226]}
// DFT_SIGNAL {random_number[227]}
// DFT_SIGNAL {random_number[228]}
// DFT_SIGNAL {random_number[229]}
// DFT_SIGNAL {random_number[230]}
// DFT_SIGNAL {random_number[231]}
// DFT_SIGNAL {random_number[232]}
// DFT_SIGNAL {random_number[233]}
// DFT_SIGNAL {random_number[234]}
// DFT_SIGNAL {random_number[235]}
// DFT_SIGNAL {random_number[236]}
// DFT_SIGNAL {random_number[237]}
// DFT_SIGNAL {random_number[238]}
// DFT_SIGNAL {random_number[239]}
// DFT_SIGNAL {random_number[240]}
// DFT_SIGNAL {random_number[241]}
// DFT_SIGNAL {random_number[242]}
// DFT_SIGNAL {random_number[243]}
// DFT_SIGNAL {random_number[244]}
// DFT_SIGNAL {random_number[245]}
// DFT_SIGNAL {random_number[246]}
// DFT_SIGNAL {random_number[247]}
// DFT_SIGNAL {random_number[248]}
// DFT_SIGNAL {random_number[249]}
// DFT_SIGNAL {random_number[250]}
// DFT_SIGNAL {random_number[251]}
// DFT_SIGNAL {random_number[252]}
// DFT_SIGNAL {random_number[253]}
// DFT_SIGNAL {random_number[254]}
// DFT_SIGNAL {random_number[255]}
// DFT_SIGNAL {clk_trng}
// DFT_SIGNAL {enable}
// DFT_SIGNAL {ready}
// DFT_SIGNAL {bist}
// DFT_SIGNAL {run}
// DFT_SIGNAL {ro_clk}

endmodule

